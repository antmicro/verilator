// Status: STUB

class uvm_report_object extends uvm_object;
endclass
