// Copyright 2023 by Antmicro Ltd.
// SPDX-License-Identifier: Apache-2.0

// Status: STUB

class uvm_report_object extends uvm_object;
endclass
