// Status: STUB

`include "base/uvm_object.svh"

class uvm_report_object extends uvm_object;
endclass
